module bo_mul_floatingpoint (
    input         clk,
    input         reset,
    input         start,
    input  [31:0] A,
    input  [31:0] B,
    output [31:0] result,
    output        overflow_flag
);

    // === T�n hi?u k?t n?i n?i b? ===
    wire MLB_significand_mult;
    wire MLB_exponent_inc;
    wire mux_en_reg;
    wire enable_reg;
    wire inc_shift_en;
    wire mux_en_rounding;
    wire enable_rounding;
    wire no_start;
    // === K?t n?i module nh�n s? th?c ===
    datapath_floatingpoint_mul mul_inst (
        .clk(clk),
        .reset(reset),
        .A(A),
        .B(B),
        .inc_shift_en(inc_shift_en),            // T�n hi?u ?i?u khi?n shift v� t?ng exp
        .mux_en_rounding(mux_en_rounding),      // Ch?n gi?a k?t qu? l�m tr�n ho?c 
        .enable_rounding(enable_rounding),
        .mux_en_reg(mux_en_reg),
        .enable_reg(enable_reg),
        .no_start(no_start),
        .MLB_exp_inc(MLB_exponent_inc),         // B�o tr�n exponent
        .MLB_significand_mult(MLB_significand_mult), // B�o c?n shift
        .result(result),
        .overflow_flag(overflow_flag)                         // K?t qu? IEEE 754
    );

    // === K?t n?i b? ?i?u khi?n ===
    control_floatingpoint_mul ctrl_inst (
        .clk(clk),
        .reset(reset),
        .start(start),
        .MLB_significand_mult(MLB_significand_mult),
        .MLB_exponent_inc(MLB_exponent_inc),
        .inc_shift_en(inc_shift_en),
        .mux_en_rounding(mux_en_rounding),
        .mux_en_reg(mux_en_reg), 
        .enable_reg(enable_reg),
        .enable_rounding(enable_rounding),
        .no_start(no_start)
    );

endmodule


